USE ieee.std_logic_1164.all;