LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

entity sad_bo is
	port (
		
	);
end sad_bo;

							
					